magic
tech scmos
timestamp 1664648421
<< nwell >>
rect -12 -5 26 29
<< polysilicon >>
rect -3 19 -1 21
rect 13 19 15 21
rect -3 -19 -1 -3
rect 13 -19 15 -3
rect -3 -37 -1 -35
rect 13 -37 15 -35
<< ndiffusion >>
rect -10 -27 -3 -19
rect -10 -31 -8 -27
rect -4 -31 -3 -27
rect -10 -35 -3 -31
rect -1 -35 13 -19
rect 15 -27 24 -19
rect 15 -31 18 -27
rect 22 -31 24 -27
rect 15 -35 24 -31
rect 18 -39 22 -35
<< pdiffusion >>
rect -10 11 -3 19
rect -10 7 -8 11
rect -4 7 -3 11
rect -10 -3 -3 7
rect -1 11 13 19
rect -1 7 4 11
rect 8 7 13 11
rect -1 -3 13 7
rect 15 11 24 19
rect 15 7 18 11
rect 22 7 24 11
rect 15 -3 24 7
<< metal1 >>
rect -18 33 33 37
rect 4 27 8 33
rect 4 11 8 23
rect -8 -15 -4 7
rect 18 -15 22 7
rect -8 -19 22 -15
rect -8 -27 -4 -19
rect 18 -39 22 -31
rect -18 -43 18 -39
rect 22 -43 33 -39
<< ntransistor >>
rect -3 -35 -1 -19
rect 13 -35 15 -19
<< ptransistor >>
rect -3 -3 -1 19
rect 13 -3 15 19
<< polycontact >>
rect -1 -11 3 -7
rect 9 -11 13 -7
<< ndcontact >>
rect -8 -31 -4 -27
rect 18 -31 22 -27
<< pdcontact >>
rect -8 7 -4 11
rect 4 7 8 11
rect 18 7 22 11
<< psubstratepcontact >>
rect 18 -43 22 -39
<< nsubstratencontact >>
rect 4 23 8 27
<< labels >>
rlabel metal1 -6 -12 -6 -12 1 out
rlabel polycontact 1 -9 1 -9 1 A
rlabel polycontact 11 -9 11 -9 1 B
rlabel metal1 13 35 13 35 5 VDD
rlabel metal1 -4 -42 -4 -42 1 GND
<< end >>
